module top
(
	input wire clk,
	input wire start,
	output wire [7:0] data
);

endmodule